entity WaitForTB is
end entity;

architecture sim of WaitForTB is
begin

    process is
    begin

        report "Boo";

    end process;

end architecture;
