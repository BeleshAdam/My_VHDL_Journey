entity t1 is
end entity;

architecture sim of t1 is
begin

    process is
    begin

        report "Hello world!";
        wait;

    end process;

end architecture;
