entity t1 is
end entity;

architecture sim of t1 is
begin

    process is
    begin




    end process;
end architecture;
